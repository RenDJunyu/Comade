    .lib './l40lp_mm_v1121.lib' tt
    .option post
    .options post_version = 9601
    .param input_rise_time=4.693E-10
    

    
    .SUBCKT PM_BUFLERMX16_DMY%I 3 7 11 15 19 23 77 79 81 83 85 87 113 GND 
C0 113 GND 0.0511389F
C1 109 GND 0.145748F
C2 100 GND 0.00706604F
C3 93 GND 0.0295604F
C4 87 GND 0.0985693F
C5 85 GND 0.0899129F
C6 83 GND 0.08989F
C7 81 GND 0.0778502F
C8 79 GND 0.0776991F
C9 77 GND 0.0986801F
C10 76 GND 0.0117316F
C11 73 GND 0.00232271F
C12 70 GND 0.00231398F
C13 67 GND 0.00147563F
C14 64 GND 0.00387201F
C15 61 GND 0.00711314F
C16 56 GND 0.0355692F
C17 50 GND 0.0324623F
C18 44 GND 0.0375109F
C19 38 GND 0.0279864F
C20 31 GND 0.0321152F
C21 23 GND 0.0684458F
C22 19 GND 0.0577454F
C23 15 GND 0.0597817F
C24 11 GND 0.0686675F
C25 7 GND 0.0675158F
C26 3 GND 0.0688496F
R27 110 113 0.250947
R28 108 109 24.0698
R29 107 108 24.0698
R30 106 107 24.0698
R31 105 106 24.0698
R32 104 105 24.0698
R33 103 104 24.0698
R34 102 103 24.0698
R35 101 102 24.0698
R36 93 110 48.011
R37 91 100 0.675381
R38 91 93 11.7827
R39 90 101 5.39284
R40 90 93 11.7827
R41 75 87 31
R42 75 76 14
R43 74 109 0.988938
R44 74 76 4
R45 72 85 31
R46 72 73 14
R47 71 107 0.988938
R48 71 73 4
R49 69 83 31
R50 69 70 14
R51 68 105 0.988938
R52 68 70 4
R53 66 81 31
R54 66 67 14
R55 65 103 0.988938
R56 65 67 4
R57 63 79 31
R58 63 64 14
R59 62 101 0.988938
R60 62 64 4
R61 60 77 31
R62 60 61 14
R63 59 100 5.75
R64 59 61 4
R65 56 108 1.64011
R66 55 73 0.46983
R67 55 56 8.19663
R68 54 76 0.46983
R69 54 56 8.19663
R70 50 106 1.64011
R71 49 70 0.46983
R72 49 50 8.19663
R73 48 73 0.46983
R74 48 50 8.19663
R75 44 104 1.64011
R76 43 67 0.46983
R77 43 44 8.19663
R78 42 70 0.46983
R79 42 44 8.19663
R80 38 102 1.64011
R81 37 64 0.46983
R82 37 38 8.19663
R83 36 67 0.46983
R84 36 38 8.19663
R85 31 110 48.011
R86 29 61 0.46983
R87 29 31 8.19663
R88 28 64 0.46983
R89 28 31 8.19663
R90 27 93 2.35765
R91 27 31 1.64011
R92 22 109 0.988938
R93 22 23 31.625
R94 18 107 0.988938
R95 18 19 31.625
R96 14 105 0.988938
R97 14 15 31.625
R98 10 103 0.988938
R99 10 11 28.75
R100 6 101 0.988938
R101 6 7 27.3125
R102 2 100 20.125
R103 2 3 30.1875
.ENDS

.SUBCKT PM_BUFLERMX16_DMY%N_1 7 8 12 13 17 18 22 23 27 28 32 33 56 60 64 68 72
+ 76 80 84 88 92 96 100 104 108 112 116 262 264 266 268 270 272 274 276 278 280
+ 282 284 286 288 290 293 GND 
C0 364 GND 0.0326676F
C1 362 GND 0.048061F
C2 359 GND 0.0617603F
C3 358 GND 0.297F
C4 341 GND 0.00395698F
C5 340 GND 0.003965F
C6 339 GND 0.00577051F
C7 338 GND 0.00158837F
C8 337 GND 0.00122733F
C9 336 GND 0.00121203F
C10 325 GND 0.0325317F
C11 321 GND 0.0344495F
C12 317 GND 0.0328064F
C13 313 GND 0.0297486F
C14 309 GND 0.100403F
C15 307 GND 0.0449082F
C16 303 GND 0.024778F
C17 298 GND 0.0319709F
C18 293 GND 0.0992959F
C19 290 GND 0.0904439F
C20 288 GND 0.0904439F
C21 286 GND 0.0904439F
C22 284 GND 0.0904439F
C23 282 GND 0.0904439F
C24 280 GND 0.0904439F
C25 278 GND 0.0904439F
C26 276 GND 0.0904439F
C27 274 GND 0.0904439F
C28 272 GND 0.0904439F
C29 270 GND 0.0749966F
C30 268 GND 0.0793778F
C31 266 GND 0.0775049F
C32 264 GND 0.0768487F
C33 262 GND 0.0983715F
C34 261 GND 0.00800616F
C35 258 GND 0.00249949F
C36 255 GND 0.00250607F
C37 252 GND 0.00250607F
C38 249 GND 0.00250607F
C39 246 GND 0.00250488F
C40 243 GND 0.00250488F
C41 240 GND 0.00250488F
C42 237 GND 0.00250607F
C43 234 GND 0.00250607F
C44 231 GND 0.00250607F
C45 228 GND 0.00294504F
C46 225 GND 0.00149672F
C47 222 GND 0.00123694F
C48 219 GND 0.00123695F
C49 215 GND 0.0120026F
C50 214 GND 0.0121354F
C51 211 GND 0.0348406F
C52 205 GND 0.035619F
C53 199 GND 0.0340607F
C54 193 GND 0.035619F
C55 187 GND 0.0340607F
C56 181 GND 0.035619F
C57 175 GND 0.0340607F
C58 169 GND 0.0356191F
C59 163 GND 0.0340607F
C60 157 GND 0.0356193F
C61 151 GND 0.0342251F
C62 145 GND 0.0301539F
C63 137 GND 0.0435327F
C64 131 GND 0.0252618F
C65 124 GND 0.0321256F
C66 116 GND 0.0687793F
C67 112 GND 0.0579937F
C68 108 GND 0.0580003F
C69 104 GND 0.0580003F
C70 100 GND 0.0580003F
C71 96 GND 0.0579991F
C72 92 GND 0.0579991F
C73 88 GND 0.0579991F
C74 84 GND 0.0577597F
C75 80 GND 0.0577011F
C76 76 GND 0.059757F
C77 72 GND 0.0658873F
C78 68 GND 0.0681717F
C79 64 GND 0.0681218F
C80 60 GND 0.068451F
C81 56 GND 0.0688677F
C82 53 GND 0.0107935F
C83 50 GND 0.0288609F
C84 49 GND 0.0148002F
C85 47 GND 0.0329456F
C86 46 GND 0.00299654F
C87 44 GND 0.00457028F
C88 43 GND 0.0120711F
C89 39 GND 0.0298717F
C90 32 GND 0.0681788F
C91 27 GND 0.0787178F
C92 22 GND 0.0696148F
C93 17 GND 0.104305F
C94 12 GND 0.101343F
C95 11 GND 0.0457476F
C96 7 GND 0.106321F
R97 359 360 1.43929
R98 355 356 24.6429
R99 354 355 24.6429
R100 353 354 24.6429
R101 352 353 24.6429
R102 351 352 24.6429
R103 350 351 24.6429
R104 349 350 24.6429
R105 348 349 24.6429
R106 347 348 24.6429
R107 346 347 24.6429
R108 345 346 24.6429
R109 344 345 24.6429
R110 343 344 24.6429
R111 342 343 24.6429
R112 324 341 0.675381
R113 324 325 11.7827
R114 323 342 5.47619
R115 323 325 11.7827
R116 320 340 0.675381
R117 320 321 11.7827
R118 319 341 0.675381
R119 319 321 11.7827
R120 316 339 0.675381
R121 316 317 11.7827
R122 315 340 0.675381
R123 315 317 11.7827
R124 312 338 0.675381
R125 312 313 11.7827
R126 311 339 0.675381
R127 311 313 11.7827
R128 309 365 0.978784
R129 307 309 96.0219
R130 306 337 0.675381
R131 306 307 11.7827
R132 305 338 0.675381
R133 305 307 11.7827
R134 302 336 0.675381
R135 302 303 11.7827
R136 301 337 0.675381
R137 301 303 11.7827
R138 298 365 32.0073
R139 296 335 2.62662
R140 296 298 11.7827
R141 295 336 0.675381
R142 295 298 11.7827
R143 260 293 31
R144 260 261 14
R145 259 358 0.83576
R146 259 261 4
R147 257 290 31
R148 257 258 14
R149 256 356 0.83576
R150 256 258 4
R151 254 288 31
R152 254 255 14
R153 253 354 0.83576
R154 253 255 4
R155 251 286 31
R156 251 252 14
R157 250 352 0.83576
R158 250 252 4
R159 248 284 31
R160 248 249 14
R161 247 350 0.83576
R162 247 249 4
R163 245 282 31
R164 245 246 14
R165 244 348 0.83576
R166 244 246 4
R167 242 280 31
R168 242 243 14
R169 241 346 0.83576
R170 241 243 4
R171 239 278 31
R172 239 240 14
R173 238 344 0.83576
R174 238 240 4
R175 236 276 31
R176 236 237 14
R177 235 342 0.83576
R178 235 237 4
R179 233 274 31
R180 233 234 14
R181 232 341 5.75
R182 232 234 4
R183 230 272 31
R184 230 231 14
R185 229 340 5.75
R186 229 231 4
R187 227 270 31
R188 227 228 14
R189 226 339 5.75
R190 226 228 4
R191 224 268 31
R192 224 225 14
R193 223 338 5.75
R194 223 225 4
R195 221 266 31
R196 221 222 14
R197 220 337 5.75
R198 220 222 4
R199 218 264 31
R200 218 219 14
R201 217 336 5.75
R202 217 219 4
R203 215 262 31
R204 215 216 10.5268
R205 214 335 3.86869
R206 214 216 2.69126
R207 210 258 0.46983
R208 210 211 8.19663
R209 209 261 0.46983
R210 209 211 8.19663
R211 208 358 24.6429
R212 208 356 24.6429
R213 208 211 1.64011
R214 205 355 1.64011
R215 204 255 0.46983
R216 204 205 8.19663
R217 203 258 0.46983
R218 203 205 8.19663
R219 199 353 1.64011
R220 198 252 0.46983
R221 198 199 8.19663
R222 197 255 0.46983
R223 197 199 8.19663
R224 193 351 1.64011
R225 192 249 0.46983
R226 192 193 8.19663
R227 191 252 0.46983
R228 191 193 8.19663
R229 187 349 1.64011
R230 186 246 0.46983
R231 186 187 8.19663
R232 185 249 0.46983
R233 185 187 8.19663
R234 181 347 1.64011
R235 180 243 0.46983
R236 180 181 8.19663
R237 179 246 0.46983
R238 179 181 8.19663
R239 175 345 1.64011
R240 174 240 0.46983
R241 174 175 8.19663
R242 173 243 0.46983
R243 173 175 8.19663
R244 169 343 1.64011
R245 168 237 0.46983
R246 168 169 8.19663
R247 167 240 0.46983
R248 167 169 8.19663
R249 162 234 0.46983
R250 162 163 8.19663
R251 161 237 0.46983
R252 161 163 8.19663
R253 160 325 2.35765
R254 160 163 1.64011
R255 156 231 0.46983
R256 156 157 8.19663
R257 155 234 0.46983
R258 155 157 8.19663
R259 154 321 2.35765
R260 154 157 1.64011
R261 150 228 0.46983
R262 150 151 8.19663
R263 149 231 0.46983
R264 149 151 8.19663
R265 148 317 2.35765
R266 148 151 1.64011
R267 144 225 0.46983
R268 144 145 8.19663
R269 143 228 0.46983
R270 143 145 8.19663
R271 142 313 2.35765
R272 142 145 1.64011
R273 137 309 96.0219
R274 136 222 0.46983
R275 136 137 8.19663
R276 135 225 0.46983
R277 135 137 8.19663
R278 134 307 2.35765
R279 134 137 1.64011
R280 130 219 0.46983
R281 130 131 8.19663
R282 129 222 0.46983
R283 129 131 8.19663
R284 128 303 2.35765
R285 128 131 1.64011
R286 124 365 32.0073
R287 122 216 1.82722
R288 122 124 8.19663
R289 121 219 0.46983
R290 121 124 8.19663
R291 120 298 2.35765
R292 120 124 1.64011
R293 115 358 0.83576
R294 115 116 31.625
R295 111 356 0.83576
R296 111 112 31.625
R297 107 354 0.83576
R298 107 108 31.625
R299 103 352 0.83576
R300 103 104 31.625
R301 99 350 0.83576
R302 99 100 31.625
R303 95 348 0.83576
R304 95 96 31.625
R305 91 346 0.83576
R306 91 92 31.625
R307 87 344 0.83576
R308 87 88 31.625
R309 83 342 0.83576
R310 83 84 30.1875
R311 79 341 20.125
R312 79 80 30.1875
R313 75 340 20.125
R314 75 76 30.1875
R315 71 339 20.125
R316 71 72 27.3125
R317 67 338 20.125
R318 67 68 27.3125
R319 63 337 20.125
R320 63 64 27.3125
R321 59 336 20.125
R322 59 60 27.3125
R323 55 335 15.1323
R324 55 56 30.1875
R325 52 365 1.206
R326 52 53 0.0756414
R327 51 362 0.24376
R328 51 53 0.0708142
R329 50 53 0.0708142
R330 48 49 0.0451841
R331 47 53 0.0756414
R332 47 48 0.741733
R333 46 364 0.0902292
R334 45 49 0.113453
R335 45 46 0.191882
R336 44 49 0.113453
R337 43 44 0.259605
R338 39 364 0.0704788
R339 39 40 1.10714
R340 36 43 0.0948811
R341 36 359 0.077228
R342 35 36 60.0137
R343 33 35 4.97329
R344 32 35 4.77273
R345 30 360 60.0137
R346 28 30 5
R347 27 30 5.21958
R348 26 50 0.365762
R349 25 26 60.0137
R350 23 25 4.77273
R351 22 25 4.77273
R352 20 362 30.0069
R353 18 20 3.16129
R354 17 20 3.16129
R355 15 364 30.0069
R356 13 15 3.16129
R357 12 15 3.16129
R358 11 40 0.133128
R359 10 11 30.0069
R360 8 10 3.16129
R361 7 10 3.16129
.ENDS

.SUBCKT PM_BUFLERMX16_DMY%O 17 18 22 23 27 28 32 33 37 38 42 43 47 48 52 53 57
+ 58 62 63 67 68 72 73 77 78 82 83 87 88 92 93 129 GND 
C0 163 GND 0.0261111F
C1 161 GND 0.0579896F
C2 159 GND 0.0538525F
C3 157 GND 0.0538525F
C4 155 GND 0.0538525F
C5 153 GND 0.0538525F
C6 151 GND 0.0417657F
C7 149 GND 0.0267289F
C8 147 GND 0.0240626F
C9 145 GND 0.0240626F
C10 143 GND 0.0240626F
C11 141 GND 0.024097F
C12 139 GND 0.0171761F
C13 135 GND 0.0206117F
C14 132 GND 0.0108168F
C15 129 GND 0.0108168F
C16 125 GND 0.0108168F
C17 122 GND 0.0111454F
C18 115 GND 0.0915835F
C19 113 GND 0.0447571F
C20 111 GND 0.0448361F
C21 109 GND 0.0448074F
C22 107 GND 0.0447653F
C23 106 GND 0.0563214F
C24 105 GND 0.0449621F
C25 104 GND 0.0284577F
C26 99 GND 0.041392F
C27 92 GND 0.0695866F
C28 87 GND 0.0784474F
C29 82 GND 0.0691975F
C30 77 GND 0.0690099F
C31 72 GND 0.0690099F
C32 67 GND 0.0690099F
C33 62 GND 0.0701221F
C34 57 GND 0.072997F
C35 52 GND 0.102831F
C36 47 GND 0.102833F
C37 42 GND 0.102833F
C38 37 GND 0.102833F
C39 32 GND 0.102866F
C40 27 GND 0.0996551F
C41 22 GND 0.103605F
C42 21 GND 0.0449427F
C43 17 GND 0.106545F
R44 136 138 1.49107
R45 134 161 0.329598
R46 134 135 0.137512
R47 133 149 0.27889
R48 133 135 0.137512
R49 131 159 0.329598
R50 131 132 0.0708142
R51 130 147 0.27889
R52 130 132 0.0708142
R53 127 157 0.329598
R54 127 129 0.0708142
R55 126 145 0.27889
R56 126 129 0.0708142
R57 124 155 0.329598
R58 124 125 0.0708142
R59 123 143 0.27889
R60 123 125 0.0708142
R61 121 153 0.329598
R62 121 122 0.0708142
R63 120 141 0.27889
R64 120 122 0.0708142
R65 119 151 0.323825
R66 117 139 0.274006
R67 117 119 0.07086
R68 116 117 0.304855
R69 115 138 0.410422
R70 115 116 0.166638
R71 114 132 0.0679243
R72 113 135 0.0138634
R73 113 114 0.496644
R74 112 129 0.0679243
R75 111 132 0.0679243
R76 111 112 0.496644
R77 110 125 0.0679243
R78 109 129 0.0679243
R79 109 110 0.496644
R80 108 122 0.0679243
R81 107 125 0.0679243
R82 107 108 0.496644
R83 106 117 0.101028
R84 105 122 0.0679243
R85 105 106 0.496644
R86 104 163 0.524956
R87 103 116 0.090014
R88 103 104 0.197978
R89 99 163 0.130834
R90 99 100 1.06378
R91 95 139 60.0137
R92 93 95 5.2324
R93 92 95 5
R94 90 136 60.0137
R95 88 90 5
R96 87 90 5.2324
R97 85 149 60.0137
R98 83 85 4.77273
R99 82 85 4.77273
R100 80 147 60.0137
R101 78 80 4.77273
R102 77 80 4.77273
R103 75 145 60.0137
R104 73 75 4.77273
R105 72 75 4.77273
R106 70 143 60.0137
R107 68 70 4.77273
R108 67 70 4.77273
R109 65 141 60.0137
R110 63 65 5
R111 62 65 5
R112 60 138 60.0137
R113 58 60 5.52632
R114 57 60 5.52632
R115 55 161 30.0069
R116 53 55 3.16129
R117 52 55 3.16129
R118 50 159 30.0069
R119 48 50 3.16129
R120 47 50 3.16129
R121 45 157 30.0069
R122 43 45 3.16129
R123 42 45 3.16129
R124 40 155 30.0069
R125 38 40 3.16129
R126 37 40 3.16129
R127 35 153 30.0069
R128 33 35 3.16129
R129 32 35 3.16129
R130 30 151 30.0069
R131 28 30 3.16129
R132 27 30 3.16129
R133 25 163 30.0069
R134 23 25 3.16129
R135 22 25 3.16129
R136 21 100 0.133128
R137 20 21 30.0069
R138 18 20 3.16129
R139 17 20 3.16129
.ENDS


.SUBCKT BUFLERMX16 O I GND VCC VCCNW 
* 
* O	O
* I	I
XMN1_B11 N_N_1_MN1_B11_D N_I_MN1_B11_G GND GND N_11_LPRVT W=2.1E-06 L=3.9324E-09
+ AD=1.512E-14 AS=2.31E-14 PD=3.675E-07 PS=6.4E-07 SA=1.1E-07 SB=7.85871E-07
+ SCA=156.898 SCB=0.0462872 SCC=0.0140624 SGA=1.4E-07 SGB=1.4E-07 SG2A=3.2E-07
+ SG2B=3.2E-07 NRD=0 NRS=0
XMN1_B11-_2 N_N_1_MN1_B11-_2_D N_I_MN1_B11-_2_G GND GND N_11_LPRVT W=1.93561E-06
+ L=3.93544E-09 AD=1.368E-14 AS=1.77333E-14 PD=3.325E-07 PS=4.38462E-07
+ SA=2.9E-07 SB=1.76E-06 SCA=167.189 SCB=0.0459543 SCC=0.0146173 SGA=1.4E-07
+ SGB=1.4E-07 SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN1_B11-_3 N_N_1_MN1_B11-_3_D N_I_MN1_B11-_3_G GND GND N_11_LPRVT W=2.06948E-06
+ L=3.92893E-09 AD=1.4381E-14 AS=1.86667E-14 PD=3.42857E-07 PS=4.61538E-07
+ SA=4.04549E-07 SB=1.61765E-06 SCA=186.925 SCB=0.0454185 SCC=0.0148011
+ SGA=1.4E-07 SGB=1.4E-07 SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN1_B11-_4 N_N_1_MN1_B11-_4_D N_I_MN1_B11-_4_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.5819E-14 AS=1.54E-14 PD=3.77143E-07 PS=3.6E-07
+ SA=4.47328E-07 SB=1.36958E-06 SCA=175.307 SCB=0.045785 SCC=0.0142548
+ SGA=1.4E-07 SGB=1.4E-07 SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN1_B11-_5 N_N_1_MN1_B11-_5_D N_I_MN1_B11-_5_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.54E-14 PD=3.6E-07 PS=3.6E-07 SA=6.92253E-07
+ SB=1.1829E-06 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN1_B11-_6 N_N_1_MN1_B11-_6_D N_I_MN1_B11-_6_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.93088E-09 AD=1.54E-14 AS=1.55023E-14 PD=3.6E-07 PS=3.68372E-07
+ SA=8.95013E-07 SB=8.12333E-07 SCA=175.307 SCB=0.045785 SCC=0.0142548
+ SGA=1.4E-07 SGB=1.4E-07 SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11 N_O_MN2_B11_D N_N_1_MN2_B11_G GND GND N_11_LPRVT W=2.13017E-06
+ L=3.9324E-09 AD=1.5015E-14 AS=1.47977E-14 PD=3.675E-07 PS=3.51628E-07
+ SA=1.10374E-06 SB=7.48082E-07 SCA=156.898 SCB=0.0462872 SCC=0.0140624
+ SGA=1.4E-07 SGB=1.4E-07 SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_2 N_O_MN2_B11-_2_D N_N_1_MN2_B11-_2_G GND GND N_11_LPRVT W=1.96405E-06
+ L=3.92973E-09 AD=1.3585E-14 AS=1.69E-14 PD=3.325E-07 PS=4.2E-07 SA=1.37E-06
+ SB=1.76E-06 SCA=167.189 SCB=0.0459543 SCC=0.0146173 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_3 N_O_MN2_B11-_3_D N_N_1_MN2_B11-_3_G GND GND N_11_LPRVT W=1.93347E-06
+ L=3.92973E-09 AD=1.33E-14 AS=1.69E-14 PD=3.3E-07 PS=4.2E-07 SA=1.55E-06
+ SB=1.76E-06 SCA=167.189 SCB=0.0459543 SCC=0.0146173 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_4 N_O_MN2_B11-_4_D N_N_1_MN2_B11-_4_G GND GND N_11_LPRVT W=1.93347E-06
+ L=3.92973E-09 AD=1.33E-14 AS=1.69E-14 PD=3.3E-07 PS=4.2E-07 SA=1.73E-06
+ SB=1.76E-06 SCA=167.189 SCB=0.0459543 SCC=0.0146173 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_5 N_O_MN2_B11-_5_D N_N_1_MN2_B11-_5_G GND GND N_11_LPRVT W=1.96405E-06
+ L=3.92973E-09 AD=1.3585E-14 AS=1.69E-14 PD=3.325E-07 PS=4.2E-07 SA=1.76E-06
+ SB=1.76E-06 SCA=167.189 SCB=0.0459543 SCC=0.0146173 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_6 N_O_MN2_B11-_6_D N_N_1_MN2_B11-_6_G GND GND N_11_LPRVT W=2.1E-06
+ L=3.92813E-09 AD=1.5015E-14 AS=1.47E-14 PD=3.675E-07 PS=3.5E-07 SA=7.48082E-07
+ SB=1.76E-06 SCA=156.898 SCB=0.0462872 SCC=0.0140624 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_7 N_O_MN2_B11-_7_D N_N_1_MN2_B11-_7_G GND GND N_11_LPRVT W=2.1E-06
+ L=3.92813E-09 AD=1.47E-14 AS=1.47E-14 PD=3.5E-07 PS=3.5E-07 SA=1.19102E-06
+ SB=1.73E-06 SCA=156.898 SCB=0.0462872 SCC=0.0140624 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_8 N_O_MN2_B11-_8_D N_N_1_MN2_B11-_8_G GND GND N_11_LPRVT W=2.1329E-06
+ L=3.94228E-09 AD=1.47E-14 AS=1.48465E-14 PD=3.5E-07 PS=3.51628E-07
+ SA=1.39502E-06 SB=1.55E-06 SCA=156.898 SCB=0.0462872 SCC=0.0140624 SGA=1.4E-07
+ SGB=1.4E-07 SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_9 N_O_MN2_B11-_9_D N_N_1_MN2_B11-_9_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.55535E-14 PD=3.6E-07 PS=3.68372E-07
+ SA=9.78285E-07 SB=1.37E-06 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07
+ SGB=1.4E-07 SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_10 N_O_MN2_B11-_10_D N_N_1_MN2_B11-_10_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.54E-14 PD=3.6E-07 PS=3.6E-07 SA=1.32241E-06
+ SB=1.19E-06 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_11 N_O_MN2_B11-_11_D N_N_1_MN2_B11-_11_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.54E-14 PD=3.6E-07 PS=3.6E-07 SA=1.47474E-06
+ SB=1.01E-06 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_12 N_O_MN2_B11-_12_D N_N_1_MN2_B11-_12_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.54E-14 PD=3.6E-07 PS=3.6E-07 SA=1.56776E-06
+ SB=8.3E-07 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_13 N_O_MN2_B11-_13_D N_N_1_MN2_B11-_13_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.54E-14 PD=3.6E-07 PS=3.6E-07 SA=1.63241E-06
+ SB=6.5E-07 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_14 N_O_MN2_B11-_14_D N_N_1_MN2_B11-_14_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.54E-14 PD=3.6E-07 PS=3.6E-07 SA=1.6806E-06
+ SB=4.7E-07 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_15 N_O_MN2_B11-_15_D N_N_1_MN2_B11-_15_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.92732E-09 AD=1.54E-14 AS=1.54E-14 PD=3.6E-07 PS=3.6E-07 SA=1.71818E-06
+ SB=2.9E-07 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMN2_B11-_16 N_O_MN2_B11-_16_D N_N_1_MN2_B11-_16_G GND GND N_11_LPRVT W=2.2E-06
+ L=3.93088E-09 AD=1.54E-14 AS=2.42E-14 PD=3.6E-07 PS=6.6E-07 SA=1.73685E-06
+ SB=1.1E-07 SCA=175.307 SCB=0.045785 SCC=0.0142548 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.8E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP1_A11 N_N_1_MP1_A11_D N_I_MP1_A11_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.01002E-09 AD=2.17E-14 AS=3.41E-14 PD=4.5E-07 PS=8.4E-07 SA=1.1E-07
+ SB=1.76E-06 SCA=118.009 SCB=0.0402304 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP1_A11-_2 N_N_1_MP1_A11-_2_D N_I_MP1_A11-_2_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=2.9E-07
+ SB=1.76E-06 SCA=117.892 SCB=0.0402188 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP1_A11-_3 N_N_1_MP1_A11-_3_D N_I_MP1_A11-_3_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=4.7E-07
+ SB=1.76E-06 SCA=117.801 SCB=0.0402137 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP1_A11-_4 N_N_1_MP1_A11-_4_D N_I_MP1_A11-_4_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=6.5E-07
+ SB=1.76E-06 SCA=117.729 SCB=0.0402115 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP1_A11-_5 N_N_1_MP1_A11-_5_D N_I_MP1_A11-_5_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=8.3E-07
+ SB=1.76E-06 SCA=117.673 SCB=0.0402105 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP1_A11-_6 N_N_1_MP1_A11-_6_D N_I_MP1_A11-_6_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.01002E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.01E-06
+ SB=1.76E-06 SCA=117.629 SCB=0.0402101 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11 N_O_MP2_A11_D N_N_1_MP2_A11_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.01002E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.19E-06
+ SB=1.76E-06 SCA=117.595 SCB=0.0402099 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_2 N_O_MP2_A11-_2_D N_N_1_MP2_A11-_2_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.37E-06
+ SB=1.76E-06 SCA=117.569 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_3 N_O_MP2_A11-_3_D N_N_1_MP2_A11-_3_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.55E-06
+ SB=1.76E-06 SCA=117.55 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_4 N_O_MP2_A11-_4_D N_N_1_MP2_A11-_4_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.73E-06
+ SB=1.76E-06 SCA=117.538 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_5 N_O_MP2_A11-_5_D N_N_1_MP2_A11-_5_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=1.76E-06 SCA=117.531 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_6 N_O_MP2_A11-_6_D N_N_1_MP2_A11-_6_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=1.76E-06 SCA=117.53 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_7 N_O_MP2_A11-_7_D N_N_1_MP2_A11-_7_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=1.73E-06 SCA=117.535 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_8 N_O_MP2_A11-_8_D N_N_1_MP2_A11-_8_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=1.55E-06 SCA=117.545 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_9 N_O_MP2_A11-_9_D N_N_1_MP2_A11-_9_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=1.37E-06 SCA=117.562 SCB=0.0402098 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_10 N_O_MP2_A11-_10_D N_N_1_MP2_A11-_10_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=1.19E-06 SCA=117.585 SCB=0.0402099 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_11 N_O_MP2_A11-_11_D N_N_1_MP2_A11-_11_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=1.01E-06 SCA=117.617 SCB=0.04021 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_12 N_O_MP2_A11-_12_D N_N_1_MP2_A11-_12_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=8.3E-07 SCA=117.657 SCB=0.0402103 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_13 N_O_MP2_A11-_13_D N_N_1_MP2_A11-_13_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=6.5E-07 SCA=117.709 SCB=0.0402111 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_14 N_O_MP2_A11-_14_D N_N_1_MP2_A11-_14_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=4.7E-07 SCA=117.775 SCB=0.0402128 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_15 N_O_MP2_A11-_15_D N_N_1_MP2_A11-_15_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.00157E-09 AD=2.17E-14 AS=2.17E-14 PD=4.5E-07 PS=4.5E-07 SA=1.76E-06
+ SB=2.9E-07 SCA=117.859 SCB=0.0402167 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.2E-07 SG2B=3.2E-07 NRD=0 NRS=0
XMP2_A11-_16 N_O_MP2_A11-_16_D N_N_1_MP2_A11-_16_G VCC VCCNW P_11_LPRVT W=3.1E-06
+ L=4.01002E-09 AD=2.17E-14 AS=3.41E-14 PD=4.5E-07 PS=8.4E-07 SA=1.76E-06
+ SB=1.1E-07 SCA=117.967 SCB=0.0402255 SCC=0.0111136 SGA=1.4E-07 SGB=1.4E-07
+ SG2A=3.8E-07 SG2B=3.2E-07 NRD=0 NRS=0
*
* FILE: NETLIST.DIST.BUFLERMX16_DMY.PXI
* CREATED: WED DEC 17 09:18:14 2014
* 
X_PM_BUFLERMX16_DMY%I N_I_MN1_B11_G N_I_MN1_B11-_2_G N_I_MN1_B11-_3_G
+ N_I_MN1_B11-_4_G N_I_MN1_B11-_5_G N_I_MN1_B11-_6_G N_I_MP1_A11_G N_I_MP1_A11-_2_G
+ N_I_MP1_A11-_3_G N_I_MP1_A11-_4_G N_I_MP1_A11-_5_G N_I_MP1_A11-_6_G I
+ GND  PM_BUFLERMX16_DMY%I
X_PM_BUFLERMX16_DMY%N_1 N_N_1_MP1_A11-_2_D N_N_1_MP1_A11_D N_N_1_MP1_A11-_4_D
+ N_N_1_MP1_A11-_3_D N_N_1_MP1_A11-_6_D N_N_1_MP1_A11-_5_D N_N_1_MN1_B11-_6_D
+ N_N_1_MN1_B11-_5_D N_N_1_MN1_B11-_2_D N_N_1_MN1_B11_D N_N_1_MN1_B11-_4_D
+ N_N_1_MN1_B11-_3_D N_N_1_MN2_B11_G N_N_1_MN2_B11-_2_G N_N_1_MN2_B11-_3_G
+ N_N_1_MN2_B11-_4_G N_N_1_MN2_B11-_5_G N_N_1_MN2_B11-_6_G N_N_1_MN2_B11-_7_G
+ N_N_1_MN2_B11-_8_G N_N_1_MN2_B11-_9_G N_N_1_MN2_B11-_10_G N_N_1_MN2_B11-_11_G
+ N_N_1_MN2_B11-_12_G N_N_1_MN2_B11-_13_G N_N_1_MN2_B11-_14_G N_N_1_MN2_B11-_15_G
+ N_N_1_MN2_B11-_16_G N_N_1_MP2_A11_G N_N_1_MP2_A11-_2_G N_N_1_MP2_A11-_3_G
+ N_N_1_MP2_A11-_4_G N_N_1_MP2_A11-_5_G N_N_1_MP2_A11-_6_G N_N_1_MP2_A11-_7_G
+ N_N_1_MP2_A11-_8_G N_N_1_MP2_A11-_9_G N_N_1_MP2_A11-_10_G N_N_1_MP2_A11-_11_G
+ N_N_1_MP2_A11-_12_G N_N_1_MP2_A11-_13_G N_N_1_MP2_A11-_14_G N_N_1_MP2_A11-_15_G
+ N_N_1_MP2_A11-_16_G GND  PM_BUFLERMX16_DMY%N_1
X_PM_BUFLERMX16_DMY%O N_O_MP2_A11-_2_D N_O_MP2_A11_D N_O_MP2_A11-_4_D
+ N_O_MP2_A11-_3_D N_O_MP2_A11-_6_D N_O_MP2_A11-_5_D N_O_MP2_A11-_8_D
+ N_O_MP2_A11-_7_D N_O_MP2_A11-_10_D N_O_MP2_A11-_9_D N_O_MP2_A11-_12_D
+ N_O_MP2_A11-_11_D N_O_MP2_A11-_14_D N_O_MP2_A11-_13_D N_O_MP2_A11-_16_D
+ N_O_MP2_A11-_15_D N_O_MN2_B11-_4_D N_O_MN2_B11-_3_D N_O_MN2_B11-_8_D
+ N_O_MN2_B11-_7_D N_O_MN2_B11-_10_D N_O_MN2_B11-_9_D N_O_MN2_B11-_12_D
+ N_O_MN2_B11-_11_D N_O_MN2_B11-_14_D N_O_MN2_B11-_13_D N_O_MN2_B11-_16_D
+ N_O_MN2_B11-_15_D N_O_MN2_B11-_2_D N_O_MN2_B11_D N_O_MN2_B11-_6_D N_O_MN2_B11-_5_D
+ O GND  PM_BUFLERMX16_DMY%O
*
.ENDS

    .temp 25
    
    .OPTION SCALE=10
    
    X_BUFLERMX16_noise noise_out noise_in noise_gnd noise_pwr noise_pwr BUFLERMX16

